magic
tech sky130A
timestamp 1615645085
<< nwell >>
rect -2 103 107 225
<< nmos >>
rect 43 25 58 67
<< pmos >>
rect 43 129 58 181
<< ndiff >>
rect 0 51 43 67
rect 0 29 20 51
rect 37 29 43 51
rect 0 25 43 29
rect 58 63 100 67
rect 58 38 66 63
rect 83 38 100 63
rect 58 25 100 38
<< pdiff >>
rect 16 175 43 181
rect 16 135 20 175
rect 37 135 43 175
rect 16 129 43 135
rect 58 177 89 181
rect 58 134 66 177
rect 83 134 89 177
rect 58 129 89 134
<< ndiffc >>
rect 20 29 37 51
rect 66 38 83 63
<< pdiffc >>
rect 20 135 37 175
rect 66 134 83 177
<< poly >>
rect 43 181 58 194
rect 43 108 58 129
rect 19 103 58 108
rect 16 86 24 103
rect 41 86 58 103
rect 19 81 58 86
rect 43 67 58 81
rect 43 12 58 25
<< polycont >>
rect 24 86 41 103
<< locali >>
rect 20 175 37 205
rect 20 127 37 135
rect 66 177 83 185
rect 66 103 83 134
rect 16 86 24 103
rect 41 86 49 103
rect 66 86 89 103
rect 66 63 83 86
rect 20 51 37 59
rect 66 30 83 38
rect 20 22 37 29
<< viali >>
rect 20 205 37 222
rect 24 86 41 103
rect 89 86 106 103
rect 20 5 37 22
<< metal1 >>
rect 0 222 107 225
rect 0 205 20 222
rect 37 205 107 222
rect 0 200 107 205
rect 18 103 47 109
rect 18 86 24 103
rect 41 86 47 103
rect 18 80 47 86
rect 83 103 112 109
rect 83 86 89 103
rect 106 86 112 103
rect 83 80 112 86
rect 0 22 100 25
rect 0 5 20 22
rect 37 5 100 22
rect 0 0 100 5
<< labels >>
rlabel metal1 0 0 100 25 0 GND!
rlabel metal1 0 200 107 225 0 Vdd!
rlabel metal1 18 80 47 109 0 Z
rlabel metal1 83 80 112 109 0 ZB
<< end >>
