magic
tech sky130A
timestamp 1615659506
<< poly >>
rect 151 556 184 561
rect 151 539 159 556
rect 176 539 184 556
rect 151 534 184 539
rect 145 501 178 506
rect 145 484 153 501
rect 170 484 178 501
rect 145 479 178 484
rect 143 444 176 449
rect 143 427 151 444
rect 168 427 176 444
rect 143 422 176 427
rect 228 438 261 443
rect 228 421 236 438
rect 253 421 261 438
rect 228 416 261 421
rect -4 152 29 157
rect -4 135 4 152
rect 21 135 29 152
rect -4 130 29 135
<< polycont >>
rect 159 539 176 556
rect 153 484 170 501
rect 151 427 168 444
rect 236 421 253 438
rect 4 135 21 152
<< locali >>
rect 151 539 159 556
rect 176 539 184 556
rect 145 484 153 501
rect 170 484 178 501
rect 143 427 151 444
rect 168 427 176 444
rect 228 421 236 438
rect 253 421 261 438
rect -4 135 4 152
rect 21 135 29 152
rect 51 148 63 166
rect 80 148 84 166
rect 102 148 106 166
rect 123 148 135 166
rect 51 110 63 128
rect 80 110 84 128
rect 0 68 33 85
rect 0 34 75 51
rect 0 0 75 17
<< viali >>
rect 159 539 176 556
rect 153 484 170 501
rect 236 421 253 438
rect 63 148 80 166
rect 106 148 123 166
rect 63 110 80 128
<< metal1 >>
rect 152 559 155 561
rect 149 536 155 559
rect 181 559 184 561
rect 152 535 155 536
rect 181 536 186 559
rect 181 535 184 536
rect 143 501 180 504
rect 143 484 153 501
rect 170 484 180 501
rect 143 481 180 484
rect 229 441 232 443
rect 226 418 232 441
rect 258 441 261 443
rect 229 417 232 418
rect 258 418 263 441
rect 258 417 261 418
rect 129 189 132 215
rect 158 189 161 215
rect 175 189 178 215
rect 204 189 207 215
rect 49 166 86 169
rect 49 148 63 166
rect 80 148 86 166
rect 49 145 86 148
rect 100 166 137 169
rect 100 148 106 166
rect 123 148 137 166
rect 100 145 137 148
rect 49 128 86 131
rect 49 110 63 128
rect 80 110 86 128
rect 100 112 160 126
rect 49 107 86 110
rect 100 28 198 42
<< rmetal1 >>
rect 100 84 198 98
rect 100 56 198 70
rect 100 0 198 14
<< via1 >>
rect 155 556 181 561
rect 155 539 159 556
rect 159 539 176 556
rect 176 539 181 556
rect 155 535 181 539
rect 232 438 258 443
rect 232 421 236 438
rect 236 421 253 438
rect 253 421 258 438
rect 232 417 258 421
rect 132 189 158 215
rect 178 189 204 215
<< metal2 >>
rect 155 561 181 564
rect 149 536 155 559
rect 181 536 186 559
rect 155 532 181 535
rect 230 444 258 449
rect 226 418 230 441
rect 258 418 263 441
rect 230 411 258 416
rect 189 341 217 346
rect 189 308 217 313
rect 257 341 285 346
rect 257 308 285 313
rect 257 273 285 278
rect 257 240 285 245
rect 132 215 158 218
rect 132 186 158 189
rect 178 215 204 218
rect 178 186 204 189
rect 184 112 198 172
rect 100 0 114 98
rect 128 0 142 98
rect 156 0 170 98
rect 184 0 198 98
<< via2 >>
rect 230 443 258 444
rect 230 417 232 443
rect 232 417 258 443
rect 230 416 258 417
rect 189 313 217 341
rect 257 313 285 341
rect 257 245 285 273
<< metal3 >>
rect 213 444 284 447
rect 213 416 230 444
rect 258 416 284 444
rect 213 413 284 416
rect 151 341 222 346
rect 151 313 189 341
rect 217 313 222 341
rect 151 308 222 313
rect 252 341 323 346
rect 252 313 257 341
rect 285 313 323 341
rect 252 308 323 313
rect 369 308 372 340
rect 404 308 444 340
rect 142 244 222 274
rect 252 273 323 278
rect 252 245 257 273
rect 285 245 323 273
rect 252 240 323 245
rect 250 180 330 210
rect 250 120 400 150
rect 250 60 400 90
rect 250 0 400 30
<< via3 >>
rect 372 308 404 340
<< metal4 >>
rect 369 340 405 377
rect 369 308 372 340
rect 404 308 405 340
rect 369 304 405 308
rect 370 180 400 260
rect 250 0 280 150
rect 310 0 340 150
rect 370 0 400 150
<< via4 >>
rect 474 440 592 558
<< metal5 >>
rect 453 558 613 570
rect 453 440 474 558
rect 592 440 613 558
rect 453 320 613 440
rect 450 0 700 160
rect 860 0 1020 250
<< end >>
